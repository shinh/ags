use std.textio.all;entity testing is end;architecture s of testing is
begin
write(output,"pong");end;